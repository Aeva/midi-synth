
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity i2s_tests is
end i2s_tests;

architecture tests of i2s_tests is
end architecture;
