

package midi is

	type frame_type is
	(
		DATA_FRAME,
		STATUS_NOTE_ON,
		STATUS_NOTE_OFF,
		STATUS_POLYPHONIC_PRESSURE,
		STATUS_CONTROL_CHANGE,
		STATUS_PROGRAM_CHANGE,
		STATUS_CHANNEL_PRESSURE,
		STATUS_PITCH_BLEND,
		STATUS_SYSTEM,
		REALTIME_TIMING_CLOCK,
		REALTIME_UNDEFINED1,
		REALTIME_START,
		REALTIME_CONTINUE,
		REALTIME_STOP,
		REALTIME_UNDEFINED2,
		REALTIME_ACTIVE_SENSE,
		REALTIME_SYSTEM_RESET
	);

	constant STATUS_OFFSET : integer := frame_type'POS(STATUS_NOTE_ON);
	constant REALTIME_OFFSET : integer := frame_type'POS(REALTIME_TIMING_CLOCK);
	
end midi;
