

package midi is

	type frame_type is
	(
		FRAME_REALTIME,
		FRAME_STATUS,
		FRAME_DATA
	);
	
	type status_message is 
	(
		STATUS_NOTE_ON,
		STATUS_NOTE_OFF,
		STATUS_POLYPHONIC_PRESSURE,
		STATUS_CONTROL_CHANGE,
		STATUS_PROGRAM_CHANGE,
		STATUS_CHANNEL_PRESSURE,
		STATUS_PITCH_BLEND,
		STATUS_SYSTEM
	);

	type realtime_message is
	(
		REALTIME_TIMING_CLOCK,
		REALTIME_UNDEFINED1,
		REALTIME_START,
		REALTIME_CONTINUE,
		REALTIME_STOP,
		REALTIME_UNDEFINED2,
		REALTIME_ACTIVE_SENSE,
		REALTIME_SYSTEM_RESET
	);	
	
end midi;
